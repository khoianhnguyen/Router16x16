`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/25/2024 10:31:34 PM
// Design Name: 
// Module Name: ROUTER
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ROUTER(
    input clk,
    input [15:0] din,
    input reset_n,
    input [15:0] frame_n,
    input [15:0] valid_n,
    output [15:0] dout,
    output [15:0] frameo_n,
    output [15:0] valido_n
    );
endmodule
