`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/03/2024 09:25:02 PM
// Design Name: 
// Module Name: Router16x16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Router16x16(
    input clk,
    input reset_n,
    input [15:0] frame_n,
    input [15:0] valid_n,
    input [15:0] din,
    output [15:0] frameo_n,
    output [15:0] valido_n,
    output [15:0] dout
    );
    wire [15:0] busy_fsm,busy_fsm1,busy_fsm2,busy_fsm3,busy_fsm4,busy_fsm5,busy_fsm6,busy_fsm7,busy_fsm8,busy_fsm9,busy_fsm10,busy_fsm11,busy_fsm12,busy_fsm13,busy_fsm14,busy_fsm15;
    wire [15:0] dout_fsm,dout_fsm1,dout_fsm2,dout_fsm3,dout_fsm4,dout_fsm5,dout_fsm6,dout_fsm7,dout_fsm8,dout_fsm9,dout_fsm10,dout_fsm11,dout_fsm12,dout_fsm13,dout_fsm14,dout_fsm15;
    wire [15:0] frameo_fsm,frameo_fsm1,frameo_fsm2,frameo_fsm3,frameo_fsm4,frameo_fsm5,frameo_fsm6,frameo_fsm7,frameo_fsm8,frameo_fsm9,frameo_fsm10,frameo_fsm11,frameo_fsm12,frameo_fsm13,frameo_fsm14,frameo_fsm15;
    wire [15:0] valido_fsm,valido_fsm1,valido_fsm2,valido_fsm3,valido_fsm4,valido_fsm5,valido_fsm6,valido_fsm7,valido_fsm8,valido_fsm9,valido_fsm10,valido_fsm11,valido_fsm12,valido_fsm13,valido_fsm14,valido_fsm15;
    
    wire [15:0] busy_arbiter,busy_arbiter1,busy_arbiter2,busy_arbiter3,busy_arbiter4,busy_arbiter5,busy_arbiter6,busy_arbiter7,busy_arbiter8,busy_arbiter9,busy_arbiter10,busy_arbiter11,busy_arbiter12,busy_arbiter13,busy_arbiter14,busy_arbiter15;
    wire [15:0] frame_arbiter,frame_arbiter1,frame_arbiter2,frame_arbiter3,frame_arbiter4,frame_arbiter5,frame_arbiter6,frame_arbiter7,frame_arbiter8,frame_arbiter9,frame_arbiter10,frame_arbiter11,frame_arbiter12,frame_arbiter13,frame_arbiter14,frame_arbiter15;
    wire [15:0] valid_arbiter,valid_arbiter1,valid_arbiter2,valid_arbiter3,valid_arbiter4,valid_arbiter5,valid_arbiter6,valid_arbiter7,valid_arbiter8,valid_arbiter9,valid_arbiter10,valid_arbiter11,valid_arbiter12,valid_arbiter13,valid_arbiter14,valid_arbiter15;
    wire [15:0] din_arbiter,din_arbiter1,din_arbiter2,din_arbiter3,din_arbiter4,din_arbiter5,din_arbiter6,din_arbiter7,din_arbiter8,din_arbiter9,din_arbiter10,din_arbiter11,din_arbiter12,din_arbiter13,din_arbiter14,din_arbiter15;
    wire [15:0] din_arbiter,din_arbiter1,din_arbiter2,din_arbiter3,din_arbiter4,din_arbiter5,din_arbiter6,din_arbiter7,din_arbiter8,din_arbiter9,din_arbiter10,din_arbiter11,din_arbiter12,din_arbiter13,din_arbiter14,din_arbiter15;
    
    fsm_decode DUT(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[0]),.valid_n(valid_n[0]),.din(din[0]),.busy(busy_fsm),.frameo_n(frameo_fsm),.valido_n(valido_fsm),.dout(dout_fsm));
    fsm_decode DUT1(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[1]),.valid_n(valid_n[1]),.din(din[1]),.busy(busy_fsm1),.frameo_n(frameo_fsm1),.valido_n(valido_fsm1),.dout(dout_fsm1));
    fsm_decode DUT2(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[2]),.valid_n(valid_n[2]),.din(din[2]),.busy(busy_fsm2),.frameo_n(frameo_fsm2),.valido_n(valido_fsm2),.dout(dout_fsm2));
    fsm_decode DUT3(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[3]),.valid_n(valid_n[3]),.din(din[3]),.busy(busy_fsm3),.frameo_n(frameo_fsm3),.valido_n(valido_fsm3),.dout(dout_fsm3));
    fsm_decode DUT4(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[4]),.valid_n(valid_n[4]),.din(din[4]),.busy(busy_fsm4),.frameo_n(frameo_fsm4),.valido_n(valido_fsm4),.dout(dout_fsm4));
    fsm_decode DUT5(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[5]),.valid_n(valid_n[5]),.din(din[5]),.busy(busy_fsm5),.frameo_n(frameo_fsm5),.valido_n(valido_fsm5),.dout(dout_fsm5));
    fsm_decode DUT6(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[6]),.valid_n(valid_n[6]),.din(din[6]),.busy(busy_fsm6),.frameo_n(frameo_fsm6),.valido_n(valido_fsm6),.dout(dout_fsm6));
    fsm_decode DUT7(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[7]),.valid_n(valid_n[7]),.din(din[7]),.busy(busy_fsm7),.frameo_n(frameo_fsm7),.valido_n(valido_fsm7),.dout(dout_fsm7));
    fsm_decode DUT8(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[8]),.valid_n(valid_n[8]),.din(din[8]),.busy(busy_fsm8),.frameo_n(frameo_fsm8),.valido_n(valido_fsm8),.dout(dout_fsm8));
    fsm_decode DUT9(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[9]),.valid_n(valid_n[9]),.din(din[9]),.busy(busy_fsm9),.frameo_n(frameo_fsm9),.valido_n(valido_fsm9),.dout(dout_fsm9));
    fsm_decode DUT10(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[10]),.valid_n(valid_n[10]),.din(din[10]),.busy(busy_fsm10),.frameo_n(frameo_fsm10),.valido_n(valido_fsm10),.dout(dout_fsm10));
    fsm_decode DUT11(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[11]),.valid_n(valid_n[11]),.din(din[11]),.busy(busy_fsm11),.frameo_n(frameo_fsm11),.valido_n(valido_fsm11),.dout(dout_fsm11));
    fsm_decode DUT12(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[12]),.valid_n(valid_n[12]),.din(din[12]),.busy(busy_fsm12),.frameo_n(frameo_fsm12),.valido_n(valido_fsm12),.dout(dout_fsm12));
    fsm_decode DUT13(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[13]),.valid_n(valid_n[13]),.din(din[13]),.busy(busy_fsm13),.frameo_n(frameo_fsm13),.valido_n(valido_fsm13),.dout(dout_fsm13));
    fsm_decode DUT14(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[14]),.valid_n(valid_n[14]),.din(din[14]),.busy(busy_fsm14),.frameo_n(frameo_fsm14),.valido_n(valido_fsm14),.dout(dout_fsm14));
    fsm_decode DUT15(.clk(clk),.reset_n(reset_n),.frame_n(frame_n[15]),.valid_n(valid_n[15]),.din(din[15]),.busy(busy_fsm15),.frameo_n(frameo_fsm15),.valido_n(valido_fsm15),.dout(dout_fsm15));
    
    Arbiter_router ADUT(.reset_n(reset_n),.din(din_arbiter),.valid_n(valid_arbiter),.frame_n(frame_arbiter),.busy(busy_arbiter),.frameo_n(frameo_n[0]),.valido_n(valido_n[0]),.dout(dout[0]));
    Arbiter_router ADUT1(.reset_n(reset_n),.din(din_arbiter1),.valid_n(valid_arbiter1),.frame_n(frame_arbiter1),.busy(busy_arbiter1),.frameo_n(frameo_n[1]),.valido_n(valido_n[1]),.dout(dout[1]));
    Arbiter_router ADUT2(.reset_n(reset_n),.din(din_arbiter2),.valid_n(valid_arbiter2),.frame_n(frame_arbiter2),.busy(busy_arbiter2),.frameo_n(frameo_n[2]),.valido_n(valido_n[2]),.dout(dout[2]));
    Arbiter_router ADUT3(.reset_n(reset_n),.din(din_arbiter3),.valid_n(valid_arbiter3),.frame_n(frame_arbiter3),.busy(busy_arbiter3),.frameo_n(frameo_n[3]),.valido_n(valido_n[3]),.dout(dout[3]));
    Arbiter_router ADUT4(.reset_n(reset_n),.din(din_arbiter4),.valid_n(valid_arbiter4),.frame_n(frame_arbiter4),.busy(busy_arbiter4),.frameo_n(frameo_n[4]),.valido_n(valido_n[4]),.dout(dout[4]));
    Arbiter_router ADUT5(.reset_n(reset_n),.din(din_arbiter5),.valid_n(valid_arbiter5),.frame_n(frame_arbiter5),.busy(busy_arbiter5),.frameo_n(frameo_n[5]),.valido_n(valido_n[5]),.dout(dout[5]));
    Arbiter_router ADUT6(.reset_n(reset_n),.din(din_arbiter6),.valid_n(valid_arbiter6),.frame_n(frame_arbiter6),.busy(busy_arbiter6),.frameo_n(frameo_n[6]),.valido_n(valido_n[6]),.dout(dout[6]));
    Arbiter_router ADUT7(.reset_n(reset_n),.din(din_arbiter7),.valid_n(valid_arbiter7),.frame_n(frame_arbiter7),.busy(busy_arbiter7),.frameo_n(frameo_n[7]),.valido_n(valido_n[7]),.dout(dout[7]));
    Arbiter_router ADUT8(.reset_n(reset_n),.din(din_arbiter8),.valid_n(valid_arbiter8),.frame_n(frame_arbiter8),.busy(busy_arbiter8),.frameo_n(frameo_n[8]),.valido_n(valido_n[8]),.dout(dout[8]));
    Arbiter_router ADUT9(.reset_n(reset_n),.din(din_arbiter9),.valid_n(valid_arbiter9),.frame_n(frame_arbiter9),.busy(busy_arbiter9),.frameo_n(frameo_n[9]),.valido_n(valido_n[9]),.dout(dout[9]));
    Arbiter_router ADUT10(.reset_n(reset_n),.din(din_arbiter10),.valid_n(valid_arbiter10),.frame_n(frame_arbiter10),.busy(busy_arbiter10),.frameo_n(frameo_n[10]),.valido_n(valido_n[10]),.dout(dout[10]));
    Arbiter_router ADUT11(.reset_n(reset_n),.din(din_arbiter11),.valid_n(valid_arbiter11),.frame_n(frame_arbiter11),.busy(busy_arbiter11),.frameo_n(frameo_n[11]),.valido_n(valido_n[11]),.dout(dout[11]));
    Arbiter_router ADUT12(.reset_n(reset_n),.din(din_arbiter12),.valid_n(valid_arbiter12),.frame_n(frame_arbiter12),.busy(busy_arbiter12),.frameo_n(frameo_n[12]),.valido_n(valido_n[12]),.dout(dout[12]));
    Arbiter_router ADUT13(.reset_n(reset_n),.din(din_arbiter13),.valid_n(valid_arbiter13),.frame_n(frame_arbiter13),.busy(busy_arbiter13),.frameo_n(frameo_n[13]),.valido_n(valido_n[13]),.dout(dout[13]));
    Arbiter_router ADUT14(.reset_n(reset_n),.din(din_arbiter14),.valid_n(valid_arbiter14),.frame_n(frame_arbiter14),.busy(busy_arbiter14),.frameo_n(frameo_n[14]),.valido_n(valido_n[14]),.dout(dout[14]));
    Arbiter_router ADUT15(.reset_n(reset_n),.din(din_arbiter15),.valid_n(valid_arbiter15),.frame_n(frame_arbiter15),.busy(busy_arbiter15),.frameo_n(frameo_n[15]),.valido_n(valido_n[15]),.dout(dout[15]));
    
    assign busy_fsm= {busy_arbiter15[0],busy_arbiter14[0],busy_arbiter13[0],busy_arbiter12[0],busy_arbiter11[0],busy_arbiter10[0],busy_arbiter9[0],busy_arbiter8[0],busy_arbiter7[0],busy_arbiter6[0],busy_arbiter5[0],busy_arbiter4[0],busy_arbiter3[0],busy_arbiter2[0],busy_arbiter1[0],busy_arbiter[0]};
    assign busy_fsm1= {busy_arbiter15[1],busy_arbiter14[1],busy_arbiter13[1],busy_arbiter12[1],busy_arbiter11[1],busy_arbiter10[1],busy_arbiter9[1],busy_arbiter8[1],busy_arbiter7[1],busy_arbiter6[1],busy_arbiter5[1],busy_arbiter4[1],busy_arbiter3[1],busy_arbiter2[1],busy_arbiter1[1],busy_arbiter[1]};
    assign busy_fsm2= {busy_arbiter15[2],busy_arbiter14[2],busy_arbiter13[2],busy_arbiter12[2],busy_arbiter11[2],busy_arbiter10[2],busy_arbiter9[2],busy_arbiter8[2],busy_arbiter7[2],busy_arbiter6[2],busy_arbiter5[2],busy_arbiter4[2],busy_arbiter3[2],busy_arbiter2[2],busy_arbiter1[2],busy_arbiter[2]};
    assign busy_fsm3= {busy_arbiter15[3],busy_arbiter14[3],busy_arbiter13[3],busy_arbiter12[3],busy_arbiter11[3],busy_arbiter10[3],busy_arbiter9[3],busy_arbiter8[3],busy_arbiter7[3],busy_arbiter6[3],busy_arbiter5[3],busy_arbiter4[3],busy_arbiter3[3],busy_arbiter2[3],busy_arbiter1[3],busy_arbiter[3]};
    assign busy_fsm4= {busy_arbiter15[4],busy_arbiter14[4],busy_arbiter13[4],busy_arbiter12[4],busy_arbiter11[4],busy_arbiter10[4],busy_arbiter9[4],busy_arbiter8[4],busy_arbiter7[4],busy_arbiter6[4],busy_arbiter5[4],busy_arbiter4[4],busy_arbiter3[4],busy_arbiter2[4],busy_arbiter1[4],busy_arbiter[4]};
    assign busy_fsm5= {busy_arbiter15[5],busy_arbiter14[5],busy_arbiter13[5],busy_arbiter12[5],busy_arbiter11[5],busy_arbiter10[5],busy_arbiter9[5],busy_arbiter8[5],busy_arbiter7[5],busy_arbiter6[5],busy_arbiter5[5],busy_arbiter4[5],busy_arbiter3[5],busy_arbiter2[5],busy_arbiter1[5],busy_arbiter[5]};
    assign busy_fsm6= {busy_arbiter15[6],busy_arbiter14[6],busy_arbiter13[6],busy_arbiter12[6],busy_arbiter11[6],busy_arbiter10[6],busy_arbiter9[6],busy_arbiter8[6],busy_arbiter7[6],busy_arbiter6[6],busy_arbiter5[6],busy_arbiter4[6],busy_arbiter3[6],busy_arbiter2[6],busy_arbiter1[6],busy_arbiter[6]};
    assign busy_fsm7= {busy_arbiter15[7],busy_arbiter14[7],busy_arbiter13[7],busy_arbiter12[7],busy_arbiter11[7],busy_arbiter10[7],busy_arbiter9[7],busy_arbiter8[7],busy_arbiter7[7],busy_arbiter6[7],busy_arbiter5[7],busy_arbiter4[7],busy_arbiter3[7],busy_arbiter2[7],busy_arbiter1[7],busy_arbiter[7]};
    assign busy_fsm8= {busy_arbiter15[8],busy_arbiter14[8],busy_arbiter13[8],busy_arbiter12[8],busy_arbiter11[8],busy_arbiter10[8],busy_arbiter9[8],busy_arbiter8[8],busy_arbiter7[8],busy_arbiter6[8],busy_arbiter5[8],busy_arbiter4[8],busy_arbiter3[8],busy_arbiter2[8],busy_arbiter1[8],busy_arbiter[8]};
    assign busy_fsm9= {busy_arbiter15[9],busy_arbiter14[9],busy_arbiter13[9],busy_arbiter12[9],busy_arbiter11[9],busy_arbiter10[9],busy_arbiter9[9],busy_arbiter8[9],busy_arbiter7[9],busy_arbiter6[9],busy_arbiter5[9],busy_arbiter4[9],busy_arbiter3[9],busy_arbiter2[9],busy_arbiter1[9],busy_arbiter[9]};
    assign busy_fsm10= {busy_arbiter15[10],busy_arbiter14[10],busy_arbiter13[10],busy_arbiter12[10],busy_arbiter11[10],busy_arbiter10[10],busy_arbiter9[10],busy_arbiter8[10],busy_arbiter7[10],busy_arbiter6[10],busy_arbiter5[10],busy_arbiter4[10],busy_arbiter3[10],busy_arbiter2[10],busy_arbiter1[10],busy_arbiter[10]};
    assign busy_fsm11= {busy_arbiter15[11],busy_arbiter14[11],busy_arbiter13[11],busy_arbiter12[11],busy_arbiter11[11],busy_arbiter10[11],busy_arbiter9[11],busy_arbiter8[11],busy_arbiter7[11],busy_arbiter6[11],busy_arbiter5[11],busy_arbiter4[11],busy_arbiter3[11],busy_arbiter2[11],busy_arbiter1[11],busy_arbiter[11]};
    assign busy_fsm12= {busy_arbiter15[12],busy_arbiter14[12],busy_arbiter13[12],busy_arbiter12[12],busy_arbiter11[12],busy_arbiter10[12],busy_arbiter9[12],busy_arbiter8[12],busy_arbiter7[12],busy_arbiter6[12],busy_arbiter5[12],busy_arbiter4[12],busy_arbiter3[12],busy_arbiter2[12],busy_arbiter1[12],busy_arbiter[12]};
    assign busy_fsm13= {busy_arbiter15[13],busy_arbiter14[13],busy_arbiter13[13],busy_arbiter12[13],busy_arbiter11[13],busy_arbiter10[13],busy_arbiter9[13],busy_arbiter8[13],busy_arbiter7[13],busy_arbiter6[13],busy_arbiter5[13],busy_arbiter4[13],busy_arbiter3[13],busy_arbiter2[13],busy_arbiter1[13],busy_arbiter[13]};
    assign busy_fsm14= {busy_arbiter15[14],busy_arbiter14[14],busy_arbiter13[14],busy_arbiter12[14],busy_arbiter11[14],busy_arbiter10[14],busy_arbiter9[14],busy_arbiter8[14],busy_arbiter7[14],busy_arbiter6[14],busy_arbiter5[14],busy_arbiter4[14],busy_arbiter3[14],busy_arbiter2[14],busy_arbiter1[14],busy_arbiter[14]};
    assign busy_fsm15= {busy_arbiter15[15],busy_arbiter14[15],busy_arbiter13[15],busy_arbiter12[15],busy_arbiter11[15],busy_arbiter10[15],busy_arbiter9[15],busy_arbiter8[15],busy_arbiter7[15],busy_arbiter6[15],busy_arbiter5[15],busy_arbiter4[15],busy_arbiter3[15],busy_arbiter2[15],busy_arbiter1[15],busy_arbiter[15]};
    
    
    
    assign din_arbiter= {dout_fsm15[0],dout_fsm14[0],dout_fsm13[0],dout_fsm12[0],dout_fsm11[0],dout_fsm10[0],dout_fsm9[0],dout_fsm8[0],dout_fsm7[0],dout_fsm6[0],dout_fsm5[0],dout_fsm4[0],dout_fsm3[0],dout_fsm2[0],dout_fsm1[0],dout_fsm[0]};
    assign din_arbiter1= {dout_fsm15[1],dout_fsm14[1],dout_fsm13[1],dout_fsm12[1],dout_fsm11[1],dout_fsm10[1],dout_fsm9[1],dout_fsm8[1],dout_fsm7[1],dout_fsm6[1],dout_fsm5[1],dout_fsm4[1],dout_fsm3[1],dout_fsm2[1],dout_fsm1[1],dout_fsm[1]};
    assign din_arbiter2= {dout_fsm15[2],dout_fsm14[2],dout_fsm13[2],dout_fsm12[2],dout_fsm11[2],dout_fsm10[2],dout_fsm9[2],dout_fsm8[2],dout_fsm7[2],dout_fsm6[2],dout_fsm5[2],dout_fsm4[2],dout_fsm3[2],dout_fsm2[2],dout_fsm1[2],dout_fsm[2]};
    assign din_arbiter3= {dout_fsm15[3],dout_fsm14[3],dout_fsm13[3],dout_fsm12[3],dout_fsm11[3],dout_fsm10[3],dout_fsm9[3],dout_fsm8[3],dout_fsm7[3],dout_fsm6[3],dout_fsm5[3],dout_fsm4[3],dout_fsm3[3],dout_fsm2[3],dout_fsm1[3],dout_fsm[3]};
    assign din_arbiter4= {dout_fsm15[4],dout_fsm14[4],dout_fsm13[4],dout_fsm12[4],dout_fsm11[4],dout_fsm10[4],dout_fsm9[4],dout_fsm8[4],dout_fsm7[4],dout_fsm6[4],dout_fsm5[4],dout_fsm4[4],dout_fsm3[4],dout_fsm2[4],dout_fsm1[4],dout_fsm[4]};
    assign din_arbiter5= {dout_fsm15[5],dout_fsm14[5],dout_fsm13[5],dout_fsm12[5],dout_fsm11[5],dout_fsm10[5],dout_fsm9[5],dout_fsm8[5],dout_fsm7[5],dout_fsm6[5],dout_fsm5[5],dout_fsm4[5],dout_fsm3[5],dout_fsm2[5],dout_fsm1[5],dout_fsm[5]};
    assign din_arbiter6= {dout_fsm15[6],dout_fsm14[6],dout_fsm13[6],dout_fsm12[6],dout_fsm11[6],dout_fsm10[6],dout_fsm9[6],dout_fsm8[6],dout_fsm7[6],dout_fsm6[6],dout_fsm5[6],dout_fsm4[6],dout_fsm3[6],dout_fsm2[6],dout_fsm1[6],dout_fsm[6]};
    assign din_arbiter7= {dout_fsm15[7],dout_fsm14[7],dout_fsm13[7],dout_fsm12[7],dout_fsm11[7],dout_fsm10[7],dout_fsm9[7],dout_fsm8[7],dout_fsm7[7],dout_fsm6[7],dout_fsm5[7],dout_fsm4[7],dout_fsm3[7],dout_fsm2[7],dout_fsm1[7],dout_fsm[7]};
    assign din_arbiter8= {dout_fsm15[8],dout_fsm14[8],dout_fsm13[8],dout_fsm12[8],dout_fsm11[8],dout_fsm10[8],dout_fsm9[8],dout_fsm8[8],dout_fsm7[8],dout_fsm6[8],dout_fsm5[8],dout_fsm4[8],dout_fsm3[8],dout_fsm2[8],dout_fsm1[8],dout_fsm[8]};
    assign din_arbiter9= {dout_fsm15[9],dout_fsm14[9],dout_fsm13[9],dout_fsm12[9],dout_fsm11[9],dout_fsm10[9],dout_fsm9[9],dout_fsm8[9],dout_fsm7[9],dout_fsm6[9],dout_fsm5[9],dout_fsm4[9],dout_fsm3[9],dout_fsm2[9],dout_fsm1[9],dout_fsm[9]};
    assign din_arbiter10= {dout_fsm15[10],dout_fsm14[10],dout_fsm13[10],dout_fsm12[10],dout_fsm11[10],dout_fsm10[10],dout_fsm9[10],dout_fsm8[10],dout_fsm7[10],dout_fsm6[10],dout_fsm5[10],dout_fsm4[10],dout_fsm3[10],dout_fsm2[10],dout_fsm1[10],dout_fsm[10]};
    assign din_arbiter11= {dout_fsm15[11],dout_fsm14[11],dout_fsm13[11],dout_fsm12[11],dout_fsm11[11],dout_fsm10[11],dout_fsm9[11],dout_fsm8[11],dout_fsm7[11],dout_fsm6[11],dout_fsm5[11],dout_fsm4[11],dout_fsm3[11],dout_fsm2[11],dout_fsm1[11],dout_fsm[11]};
    assign din_arbiter12= {dout_fsm15[12],dout_fsm14[12],dout_fsm13[12],dout_fsm12[12],dout_fsm11[12],dout_fsm10[12],dout_fsm9[12],dout_fsm8[12],dout_fsm7[12],dout_fsm6[12],dout_fsm5[12],dout_fsm4[12],dout_fsm3[12],dout_fsm2[12],dout_fsm1[12],dout_fsm[12]};
    assign din_arbiter13= {dout_fsm15[13],dout_fsm14[13],dout_fsm13[13],dout_fsm12[13],dout_fsm11[13],dout_fsm10[13],dout_fsm9[13],dout_fsm8[13],dout_fsm7[13],dout_fsm6[13],dout_fsm5[13],dout_fsm4[13],dout_fsm3[13],dout_fsm2[13],dout_fsm1[13],dout_fsm[13]};
    assign din_arbiter14= {dout_fsm15[14],dout_fsm14[14],dout_fsm13[14],dout_fsm12[14],dout_fsm11[14],dout_fsm10[14],dout_fsm9[14],dout_fsm8[14],dout_fsm7[14],dout_fsm6[14],dout_fsm5[14],dout_fsm4[14],dout_fsm3[14],dout_fsm2[14],dout_fsm1[14],dout_fsm[14]};
    assign din_arbiter15= {dout_fsm15[15],dout_fsm14[15],dout_fsm13[15],dout_fsm12[15],dout_fsm11[15],dout_fsm10[15],dout_fsm9[15],dout_fsm8[15],dout_fsm7[15],dout_fsm6[15],dout_fsm5[15],dout_fsm4[15],dout_fsm3[15],dout_fsm2[15],dout_fsm1[15],dout_fsm[15]};
    
     
    assign valid_arbiter= {valido_fsm15[0],valido_fsm14[0],valido_fsm13[0],valido_fsm12[0],valido_fsm11[0],valido_fsm10[0],valido_fsm9[0],valido_fsm8[0],valido_fsm7[0],valido_fsm6[0],valido_fsm5[0],valido_fsm4[0],valido_fsm3[0],valido_fsm2[0],valido_fsm1[0],valido_fsm[0]};
    assign valid_arbiter1= {valido_fsm15[1],valido_fsm14[1],valido_fsm13[1],valido_fsm12[1],valido_fsm11[1],valido_fsm10[1],valido_fsm9[1],valido_fsm8[1],valido_fsm7[1],valido_fsm6[1],valido_fsm5[1],valido_fsm4[1],valido_fsm3[1],valido_fsm2[1],valido_fsm1[1],valido_fsm[1]};
    assign valid_arbiter2= {valido_fsm15[2],valido_fsm14[2],valido_fsm13[2],valido_fsm12[2],valido_fsm11[2],valido_fsm10[2],valido_fsm9[2],valido_fsm8[2],valido_fsm7[2],valido_fsm6[2],valido_fsm5[2],valido_fsm4[2],valido_fsm3[2],valido_fsm2[2],valido_fsm1[2],valido_fsm[2]};
    assign valid_arbiter3= {valido_fsm15[3],valido_fsm14[3],valido_fsm13[3],valido_fsm12[3],valido_fsm11[3],valido_fsm10[3],valido_fsm9[3],valido_fsm8[3],valido_fsm7[3],valido_fsm6[3],valido_fsm5[3],valido_fsm4[3],valido_fsm3[3],valido_fsm2[3],valido_fsm1[3],valido_fsm[3]};
    assign valid_arbiter4= {valido_fsm15[4],valido_fsm14[4],valido_fsm13[4],valido_fsm12[4],valido_fsm11[4],valido_fsm10[4],valido_fsm9[4],valido_fsm8[4],valido_fsm7[4],valido_fsm6[4],valido_fsm5[4],valido_fsm4[4],valido_fsm3[4],valido_fsm2[4],valido_fsm1[4],valido_fsm[4]};
    assign valid_arbiter5= {valido_fsm15[5],valido_fsm14[5],valido_fsm13[5],valido_fsm12[5],valido_fsm11[5],valido_fsm10[5],valido_fsm9[5],valido_fsm8[5],valido_fsm7[5],valido_fsm6[5],valido_fsm5[5],valido_fsm4[5],valido_fsm3[5],valido_fsm2[5],valido_fsm1[5],valido_fsm[5]};
    assign valid_arbiter6= {valido_fsm15[6],valido_fsm14[6],valido_fsm13[6],valido_fsm12[6],valido_fsm11[6],valido_fsm10[6],valido_fsm9[6],valido_fsm8[6],valido_fsm7[6],valido_fsm6[6],valido_fsm5[6],valido_fsm4[6],valido_fsm3[6],valido_fsm2[6],valido_fsm1[6],valido_fsm[6]};
    assign valid_arbiter7= {valido_fsm15[7],valido_fsm14[7],valido_fsm13[7],valido_fsm12[7],valido_fsm11[7],valido_fsm10[7],valido_fsm9[7],valido_fsm8[7],valido_fsm7[7],valido_fsm6[7],valido_fsm5[7],valido_fsm4[7],valido_fsm3[7],valido_fsm2[7],valido_fsm1[7],valido_fsm[7]};
    assign valid_arbiter8= {valido_fsm15[8],valido_fsm14[8],valido_fsm13[8],valido_fsm12[8],valido_fsm11[8],valido_fsm10[8],valido_fsm9[8],valido_fsm8[8],valido_fsm7[8],valido_fsm6[8],valido_fsm5[8],valido_fsm4[8],valido_fsm3[8],valido_fsm2[8],valido_fsm1[8],valido_fsm[8]};
    assign valid_arbiter9= {valido_fsm15[9],valido_fsm14[9],valido_fsm13[9],valido_fsm12[9],valido_fsm11[9],valido_fsm10[9],valido_fsm9[9],valido_fsm8[9],valido_fsm7[9],valido_fsm6[9],valido_fsm5[9],valido_fsm4[9],valido_fsm3[9],valido_fsm2[9],valido_fsm1[9],valido_fsm[9]};
    assign valid_arbiter10= {valido_fsm15[10],valido_fsm14[10],valido_fsm13[10],valido_fsm12[10],valido_fsm11[10],valido_fsm10[10],valido_fsm9[10],valido_fsm8[10],valido_fsm7[10],valido_fsm6[10],valido_fsm5[10],valido_fsm4[10],valido_fsm3[10],valido_fsm2[10],valido_fsm1[10],valido_fsm[10]};
    assign valid_arbiter11= {valido_fsm15[11],valido_fsm14[11],valido_fsm13[11],valido_fsm12[11],valido_fsm11[11],valido_fsm10[11],valido_fsm9[11],valido_fsm8[11],valido_fsm7[11],valido_fsm6[11],valido_fsm5[11],valido_fsm4[11],valido_fsm3[11],valido_fsm2[11],valido_fsm1[11],valido_fsm[11]};
    assign valid_arbiter12= {valido_fsm15[12],valido_fsm14[12],valido_fsm13[12],valido_fsm12[12],valido_fsm11[12],valido_fsm10[12],valido_fsm9[12],valido_fsm8[12],valido_fsm7[12],valido_fsm6[12],valido_fsm5[12],valido_fsm4[12],valido_fsm3[12],valido_fsm2[12],valido_fsm1[12],valido_fsm[12]};
    assign valid_arbiter13= {valido_fsm15[13],valido_fsm14[13],valido_fsm13[13],valido_fsm12[13],valido_fsm11[13],valido_fsm10[13],valido_fsm9[13],valido_fsm8[13],valido_fsm7[13],valido_fsm6[13],valido_fsm5[13],valido_fsm4[13],valido_fsm3[13],valido_fsm2[13],valido_fsm1[13],valido_fsm[13]};
    assign valid_arbiter14= {valido_fsm15[14],valido_fsm14[14],valido_fsm13[14],valido_fsm12[14],valido_fsm11[14],valido_fsm10[14],valido_fsm9[14],valido_fsm8[14],valido_fsm7[14],valido_fsm6[14],valido_fsm5[14],valido_fsm4[14],valido_fsm3[14],valido_fsm2[14],valido_fsm1[14],valido_fsm[14]};
    assign valid_arbiter15= {valido_fsm15[15],valido_fsm14[15],valido_fsm13[15],valido_fsm12[15],valido_fsm11[15],valido_fsm10[15],valido_fsm9[15],valido_fsm8[15],valido_fsm7[15],valido_fsm6[15],valido_fsm5[15],valido_fsm4[15],valido_fsm3[15],valido_fsm2[15],valido_fsm1[15],valido_fsm[15]};
   
   
    assign frame_arbiter= {frameo_fsm15[0],frameo_fsm14[0],frameo_fsm13[0],frameo_fsm12[0],frameo_fsm11[0],frameo_fsm10[0],frameo_fsm9[0],frameo_fsm8[0],frameo_fsm7[0],frameo_fsm6[0],frameo_fsm5[0],frameo_fsm4[0],frameo_fsm3[0],frameo_fsm2[0],frameo_fsm1[0],frameo_fsm[0]};
    assign frame_arbiter1= {frameo_fsm15[1],frameo_fsm14[1],frameo_fsm13[1],frameo_fsm12[1],frameo_fsm11[1],frameo_fsm10[1],frameo_fsm9[1],frameo_fsm8[1],frameo_fsm7[1],frameo_fsm6[1],frameo_fsm5[1],frameo_fsm4[1],frameo_fsm3[1],frameo_fsm2[1],frameo_fsm1[1],frameo_fsm[1]};
    assign frame_arbiter2= {frameo_fsm15[2],frameo_fsm14[2],frameo_fsm13[2],frameo_fsm12[2],frameo_fsm11[2],frameo_fsm10[2],frameo_fsm9[2],frameo_fsm8[2],frameo_fsm7[2],frameo_fsm6[2],frameo_fsm5[2],frameo_fsm4[2],frameo_fsm3[2],frameo_fsm2[2],frameo_fsm1[2],frameo_fsm[2]};
    assign frame_arbiter3= {frameo_fsm15[3],frameo_fsm14[3],frameo_fsm13[3],frameo_fsm12[3],frameo_fsm11[3],frameo_fsm10[3],frameo_fsm9[3],frameo_fsm8[3],frameo_fsm7[3],frameo_fsm6[3],frameo_fsm5[3],frameo_fsm4[3],frameo_fsm3[3],frameo_fsm2[3],frameo_fsm1[3],frameo_fsm[3]};
    assign frame_arbiter4= {frameo_fsm15[4],frameo_fsm14[4],frameo_fsm13[4],frameo_fsm12[4],frameo_fsm11[4],frameo_fsm10[4],frameo_fsm9[4],frameo_fsm8[4],frameo_fsm7[4],frameo_fsm6[4],frameo_fsm5[4],frameo_fsm4[4],frameo_fsm3[4],frameo_fsm2[4],frameo_fsm1[4],frameo_fsm[4]};
    assign frame_arbiter5= {frameo_fsm15[5],frameo_fsm14[5],frameo_fsm13[5],frameo_fsm12[5],frameo_fsm11[5],frameo_fsm10[5],frameo_fsm9[5],frameo_fsm8[5],frameo_fsm7[5],frameo_fsm6[5],frameo_fsm5[5],frameo_fsm4[5],frameo_fsm3[5],frameo_fsm2[5],frameo_fsm1[5],frameo_fsm[5]};
    assign frame_arbiter6= {frameo_fsm15[6],frameo_fsm14[6],frameo_fsm13[6],frameo_fsm12[6],frameo_fsm11[6],frameo_fsm10[6],frameo_fsm9[6],frameo_fsm8[6],frameo_fsm7[6],frameo_fsm6[6],frameo_fsm5[6],frameo_fsm4[6],frameo_fsm3[6],frameo_fsm2[6],frameo_fsm1[6],frameo_fsm[6]};
    assign frame_arbiter7= {frameo_fsm15[7],frameo_fsm14[7],frameo_fsm13[7],frameo_fsm12[7],frameo_fsm11[7],frameo_fsm10[7],frameo_fsm9[7],frameo_fsm8[7],frameo_fsm7[7],frameo_fsm6[7],frameo_fsm5[7],frameo_fsm4[7],frameo_fsm3[7],frameo_fsm2[7],frameo_fsm1[7],frameo_fsm[7]};
    assign frame_arbiter8= {frameo_fsm15[8],frameo_fsm14[8],frameo_fsm13[8],frameo_fsm12[8],frameo_fsm11[8],frameo_fsm10[8],frameo_fsm9[8],frameo_fsm8[8],frameo_fsm7[8],frameo_fsm6[8],frameo_fsm5[8],frameo_fsm4[8],frameo_fsm3[8],frameo_fsm2[8],frameo_fsm1[8],frameo_fsm[8]};
    assign frame_arbiter9= {frameo_fsm15[9],frameo_fsm14[9],frameo_fsm13[9],frameo_fsm12[9],frameo_fsm11[9],frameo_fsm10[9],frameo_fsm9[9],frameo_fsm8[9],frameo_fsm7[9],frameo_fsm6[9],frameo_fsm5[9],frameo_fsm4[9],frameo_fsm3[9],frameo_fsm2[9],frameo_fsm1[9],frameo_fsm[9]};
    assign frame_arbiter10= {frameo_fsm15[10],frameo_fsm14[10],frameo_fsm13[10],frameo_fsm12[10],frameo_fsm11[10],frameo_fsm10[10],frameo_fsm9[10],frameo_fsm8[10],frameo_fsm7[10],frameo_fsm6[10],frameo_fsm5[10],frameo_fsm4[10],frameo_fsm3[10],frameo_fsm2[10],frameo_fsm1[10],frameo_fsm[10]};
    assign frame_arbiter11= {frameo_fsm15[11],frameo_fsm14[11],frameo_fsm13[11],frameo_fsm12[11],frameo_fsm11[11],frameo_fsm10[11],frameo_fsm9[11],frameo_fsm8[11],frameo_fsm7[11],frameo_fsm6[11],frameo_fsm5[11],frameo_fsm4[11],frameo_fsm3[11],frameo_fsm2[11],frameo_fsm1[11],frameo_fsm[11]};
    assign frame_arbiter12= {frameo_fsm15[12],frameo_fsm14[12],frameo_fsm13[12],frameo_fsm12[12],frameo_fsm11[12],frameo_fsm10[12],frameo_fsm9[12],frameo_fsm8[12],frameo_fsm7[12],frameo_fsm6[12],frameo_fsm5[12],frameo_fsm4[12],frameo_fsm3[12],frameo_fsm2[12],frameo_fsm1[12],frameo_fsm[12]};
    assign frame_arbiter13= {frameo_fsm15[13],frameo_fsm14[13],frameo_fsm13[13],frameo_fsm12[13],frameo_fsm11[13],frameo_fsm10[13],frameo_fsm9[13],frameo_fsm8[13],frameo_fsm7[13],frameo_fsm6[13],frameo_fsm5[13],frameo_fsm4[13],frameo_fsm3[13],frameo_fsm2[13],frameo_fsm1[13],frameo_fsm[13]};
    assign frame_arbiter14= {frameo_fsm15[14],frameo_fsm14[14],frameo_fsm13[14],frameo_fsm12[14],frameo_fsm11[14],frameo_fsm10[14],frameo_fsm9[14],frameo_fsm8[14],frameo_fsm7[14],frameo_fsm6[14],frameo_fsm5[14],frameo_fsm4[14],frameo_fsm3[14],frameo_fsm2[14],frameo_fsm1[14],frameo_fsm[14]};
    assign frame_arbiter15= {frameo_fsm15[15],frameo_fsm14[15],frameo_fsm13[15],frameo_fsm12[15],frameo_fsm11[15],frameo_fsm10[15],frameo_fsm9[15],frameo_fsm8[15],frameo_fsm7[15],frameo_fsm6[15],frameo_fsm5[15],frameo_fsm4[15],frameo_fsm3[15],frameo_fsm2[15],frameo_fsm1[15],frameo_fsm[15]};
endmodule
